`include "syn_interface.sv"
`include "syn_seq_item.sv"
`include "syn_sequence.sv"
`include "syn_sequencer.sv"
`include "syn_driver.sv"
`include "syn_monitor.sv"
`include "syn_agent.sv"
`include "syn_env.sv"
`include "syn_test.sv"
